//
//    Copyright (C) 2022  Jakub Hladik
//
//    This program is free software: you can redistribute it and/or modify
//    it under the terms of the GNU General Public License as published by
//    the Free Software Foundation, either version 3 of the License, or
//    (at your option) any later version.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    You should have received a copy of the GNU General Public License
//    along with this program.  If not, see <https://www.gnu.org/licenses/>.
//

`default_nettype none

module PS7 (
    /* verilator lint_off UNUSED */
    /* verilator lint_off UNDRIVEN */
    output logic [ 1:0] DMA0DATYPE,
    output logic        DMA0DAVALID,
    output logic        DMA0DRREADY,
    output logic        DMA0RSTN,
    output logic [ 1:0] DMA1DATYPE,
    output logic        DMA1DAVALID,
    output logic        DMA1DRREADY,
    output logic        DMA1RSTN,
    output logic [ 1:0] DMA2DATYPE,
    output logic        DMA2DAVALID,
    output logic        DMA2DRREADY,
    output logic        DMA2RSTN,
    output logic [ 1:0] DMA3DATYPE,
    output logic        DMA3DAVALID,
    output logic        DMA3DRREADY,
    output logic        DMA3RSTN,
    output logic        EMIOCAN0PHYTX,
    output logic        EMIOCAN1PHYTX,
    output logic [ 7:0] EMIOENET0GMIITXD,
    output logic        EMIOENET0GMIITXEN,
    output logic        EMIOENET0GMIITXER,
    output logic        EMIOENET0MDIOMDC,
    output logic        EMIOENET0MDIOO,
    output logic        EMIOENET0MDIOTN,
    output logic        EMIOENET0PTPDELAYREQRX,
    output logic        EMIOENET0PTPDELAYREQTX,
    output logic        EMIOENET0PTPPDELAYREQRX,
    output logic        EMIOENET0PTPPDELAYREQTX,
    output logic        EMIOENET0PTPPDELAYRESPRX,
    output logic        EMIOENET0PTPPDELAYRESPTX,
    output logic        EMIOENET0PTPSYNCFRAMERX,
    output logic        EMIOENET0PTPSYNCFRAMETX,
    output logic        EMIOENET0SOFRX,
    output logic        EMIOENET0SOFTX,
    output logic [ 7:0] EMIOENET1GMIITXD,
    output logic        EMIOENET1GMIITXEN,
    output logic        EMIOENET1GMIITXER,
    output logic        EMIOENET1MDIOMDC,
    output logic        EMIOENET1MDIOO,
    output logic        EMIOENET1MDIOTN,
    output logic        EMIOENET1PTPDELAYREQRX,
    output logic        EMIOENET1PTPDELAYREQTX,
    output logic        EMIOENET1PTPPDELAYREQRX,
    output logic        EMIOENET1PTPPDELAYREQTX,
    output logic        EMIOENET1PTPPDELAYRESPRX,
    output logic        EMIOENET1PTPPDELAYRESPTX,
    output logic        EMIOENET1PTPSYNCFRAMERX,
    output logic        EMIOENET1PTPSYNCFRAMETX,
    output logic        EMIOENET1SOFRX,
    output logic        EMIOENET1SOFTX,
    output logic [63:0] EMIOGPIOO,
    output logic [63:0] EMIOGPIOTN,
    output logic        EMIOI2C0SCLO,
    output logic        EMIOI2C0SCLTN,
    output logic        EMIOI2C0SDAO,
    output logic        EMIOI2C0SDATN,
    output logic        EMIOI2C1SCLO,
    output logic        EMIOI2C1SCLTN,
    output logic        EMIOI2C1SDAO,
    output logic        EMIOI2C1SDATN,
    output logic        EMIOPJTAGTDO,
    output logic        EMIOPJTAGTDTN,
    output logic        EMIOSDIO0BUSPOW,
    output logic [ 2:0] EMIOSDIO0BUSVOLT,
    output logic        EMIOSDIO0CLK,
    output logic        EMIOSDIO0CMDO,
    output logic        EMIOSDIO0CMDTN,
    output logic [ 3:0] EMIOSDIO0DATAO,
    output logic [ 3:0] EMIOSDIO0DATATN,
    output logic        EMIOSDIO0LED,
    output logic        EMIOSDIO1BUSPOW,
    output logic [ 2:0] EMIOSDIO1BUSVOLT,
    output logic        EMIOSDIO1CLK,
    output logic        EMIOSDIO1CMDO,
    output logic        EMIOSDIO1CMDTN,
    output logic [ 3:0] EMIOSDIO1DATAO,
    output logic [ 3:0] EMIOSDIO1DATATN,
    output logic        EMIOSDIO1LED,
    output logic        EMIOSPI0MO,
    output logic        EMIOSPI0MOTN,
    output logic        EMIOSPI0SCLKO,
    output logic        EMIOSPI0SCLKTN,
    output logic        EMIOSPI0SO,
    output logic        EMIOSPI0SSNTN,
    output logic [ 2:0] EMIOSPI0SSON,
    output logic        EMIOSPI0STN,
    output logic        EMIOSPI1MO,
    output logic        EMIOSPI1MOTN,
    output logic        EMIOSPI1SCLKO,
    output logic        EMIOSPI1SCLKTN,
    output logic        EMIOSPI1SO,
    output logic        EMIOSPI1SSNTN,
    output logic [ 2:0] EMIOSPI1SSON,
    output logic        EMIOSPI1STN,
    output logic        EMIOTRACECTL,
    output logic [31:0] EMIOTRACEDATA,
    output logic [ 2:0] EMIOTTC0WAVEO,
    output logic [ 2:0] EMIOTTC1WAVEO,
    output logic        EMIOUART0DTRN,
    output logic        EMIOUART0RTSN,
    output logic        EMIOUART0TX,
    output logic        EMIOUART1DTRN,
    output logic        EMIOUART1RTSN,
    output logic        EMIOUART1TX,
    output logic [ 1:0] EMIOUSB0PORTINDCTL,
    output logic        EMIOUSB0VBUSPWRSELECT,
    output logic [ 1:0] EMIOUSB1PORTINDCTL,
    output logic        EMIOUSB1VBUSPWRSELECT,
    output logic        EMIOWDTRSTO,
    output logic        EVENTEVENTO,
    output logic [ 1:0] EVENTSTANDBYWFE,
    output logic [ 1:0] EVENTSTANDBYWFI,
    output logic [ 3:0] FCLKCLK,
    output logic [ 3:0] FCLKRESETN,
    output logic [ 3:0] FTMTF2PTRIGACK,
    output logic [31:0] FTMTP2FDEBUG,
    output logic [ 3:0] FTMTP2FTRIG,
    output logic [28:0] IRQP2F,
    output logic [31:0] MAXIGP0ARADDR,
    output logic [ 1:0] MAXIGP0ARBURST,
    output logic [ 3:0] MAXIGP0ARCACHE,
    output logic        MAXIGP0ARESETN,
    output logic [11:0] MAXIGP0ARID,
    output logic [ 3:0] MAXIGP0ARLEN,
    output logic [ 1:0] MAXIGP0ARLOCK,
    output logic [ 2:0] MAXIGP0ARPROT,
    output logic [ 3:0] MAXIGP0ARQOS,
    output logic [ 1:0] MAXIGP0ARSIZE,
    output logic        MAXIGP0ARVALID,
    output logic [31:0] MAXIGP0AWADDR,
    output logic [ 1:0] MAXIGP0AWBURST,
    output logic [ 3:0] MAXIGP0AWCACHE,
    output logic [11:0] MAXIGP0AWID,
    output logic [ 3:0] MAXIGP0AWLEN,
    output logic [ 1:0] MAXIGP0AWLOCK,
    output logic [ 2:0] MAXIGP0AWPROT,
    output logic [ 3:0] MAXIGP0AWQOS,
    output logic [ 1:0] MAXIGP0AWSIZE,
    output logic        MAXIGP0AWVALID,
    output logic        MAXIGP0BREADY,
    output logic        MAXIGP0RREADY,
    output logic [31:0] MAXIGP0WDATA,
    output logic [11:0] MAXIGP0WID,
    output logic        MAXIGP0WLAST,
    output logic [ 3:0] MAXIGP0WSTRB,
    output logic        MAXIGP0WVALID,
    output logic [31:0] MAXIGP1ARADDR,
    output logic [ 1:0] MAXIGP1ARBURST,
    output logic [ 3:0] MAXIGP1ARCACHE,
    output logic        MAXIGP1ARESETN,
    output logic [11:0] MAXIGP1ARID,
    output logic [ 3:0] MAXIGP1ARLEN,
    output logic [ 1:0] MAXIGP1ARLOCK,
    output logic [ 2:0] MAXIGP1ARPROT,
    output logic [ 3:0] MAXIGP1ARQOS,
    output logic [ 1:0] MAXIGP1ARSIZE,
    output logic        MAXIGP1ARVALID,
    output logic [31:0] MAXIGP1AWADDR,
    output logic [ 1:0] MAXIGP1AWBURST,
    output logic [ 3:0] MAXIGP1AWCACHE,
    output logic [11:0] MAXIGP1AWID,
    output logic [ 3:0] MAXIGP1AWLEN,
    output logic [ 1:0] MAXIGP1AWLOCK,
    output logic [ 2:0] MAXIGP1AWPROT,
    output logic [ 3:0] MAXIGP1AWQOS,
    output logic [ 1:0] MAXIGP1AWSIZE,
    output logic        MAXIGP1AWVALID,
    output logic        MAXIGP1BREADY,
    output logic        MAXIGP1RREADY,
    output logic [31:0] MAXIGP1WDATA,
    output logic [11:0] MAXIGP1WID,
    output logic        MAXIGP1WLAST,
    output logic [ 3:0] MAXIGP1WSTRB,
    output logic        MAXIGP1WVALID,
    output logic        SAXIACPARESETN,
    output logic        SAXIACPARREADY,
    output logic        SAXIACPAWREADY,
    output logic [ 2:0] SAXIACPBID,
    output logic [ 1:0] SAXIACPBRESP,
    output logic        SAXIACPBVALID,
    output logic [63:0] SAXIACPRDATA,
    output logic [ 2:0] SAXIACPRID,
    output logic        SAXIACPRLAST,
    output logic [ 1:0] SAXIACPRRESP,
    output logic        SAXIACPRVALID,
    output logic        SAXIACPWREADY,
    output logic        SAXIGP0ARESETN,
    output logic        SAXIGP0ARREADY,
    output logic        SAXIGP0AWREADY,
    output logic [ 5:0] SAXIGP0BID,
    output logic [ 1:0] SAXIGP0BRESP,
    output logic        SAXIGP0BVALID,
    output logic [31:0] SAXIGP0RDATA,
    output logic [ 5:0] SAXIGP0RID,
    output logic        SAXIGP0RLAST,
    output logic [ 1:0] SAXIGP0RRESP,
    output logic        SAXIGP0RVALID,
    output logic        SAXIGP0WREADY,
    output logic        SAXIGP1ARESETN,
    output logic        SAXIGP1ARREADY,
    output logic        SAXIGP1AWREADY,
    output logic [ 5:0] SAXIGP1BID,
    output logic [ 1:0] SAXIGP1BRESP,
    output logic        SAXIGP1BVALID,
    output logic [31:0] SAXIGP1RDATA,
    output logic [ 5:0] SAXIGP1RID,
    output logic        SAXIGP1RLAST,
    output logic [ 1:0] SAXIGP1RRESP,
    output logic        SAXIGP1RVALID,
    output logic        SAXIGP1WREADY,
    output logic        SAXIHP0ARESETN,
    output logic        SAXIHP0ARREADY,
    output logic        SAXIHP0AWREADY,
    output logic [ 5:0] SAXIHP0BID,
    output logic [ 1:0] SAXIHP0BRESP,
    output logic        SAXIHP0BVALID,
    output logic [ 2:0] SAXIHP0RACOUNT,
    output logic [ 7:0] SAXIHP0RCOUNT,
    output logic [63:0] SAXIHP0RDATA,
    output logic [ 5:0] SAXIHP0RID,
    output logic        SAXIHP0RLAST,
    output logic [ 1:0] SAXIHP0RRESP,
    output logic        SAXIHP0RVALID,
    output logic [ 5:0] SAXIHP0WACOUNT,
    output logic [ 7:0] SAXIHP0WCOUNT,
    output logic        SAXIHP0WREADY,
    output logic        SAXIHP1ARESETN,
    output logic        SAXIHP1ARREADY,
    output logic        SAXIHP1AWREADY,
    output logic [ 5:0] SAXIHP1BID,
    output logic [ 1:0] SAXIHP1BRESP,
    output logic        SAXIHP1BVALID,
    output logic [ 2:0] SAXIHP1RACOUNT,
    output logic [ 7:0] SAXIHP1RCOUNT,
    output logic [63:0] SAXIHP1RDATA,
    output logic [ 5:0] SAXIHP1RID,
    output logic        SAXIHP1RLAST,
    output logic [ 1:0] SAXIHP1RRESP,
    output logic        SAXIHP1RVALID,
    output logic [ 5:0] SAXIHP1WACOUNT,
    output logic [ 7:0] SAXIHP1WCOUNT,
    output logic        SAXIHP1WREADY,
    output logic        SAXIHP2ARESETN,
    output logic        SAXIHP2ARREADY,
    output logic        SAXIHP2AWREADY,
    output logic [ 5:0] SAXIHP2BID,
    output logic [ 1:0] SAXIHP2BRESP,
    output logic        SAXIHP2BVALID,
    output logic [ 2:0] SAXIHP2RACOUNT,
    output logic [ 7:0] SAXIHP2RCOUNT,
    output logic [63:0] SAXIHP2RDATA,
    output logic [ 5:0] SAXIHP2RID,
    output logic        SAXIHP2RLAST,
    output logic [ 1:0] SAXIHP2RRESP,
    output logic        SAXIHP2RVALID,
    output logic [ 5:0] SAXIHP2WACOUNT,
    output logic [ 7:0] SAXIHP2WCOUNT,
    output logic        SAXIHP2WREADY,
    output logic        SAXIHP3ARESETN,
    output logic        SAXIHP3ARREADY,
    output logic        SAXIHP3AWREADY,
    output logic [ 5:0] SAXIHP3BID,
    output logic [ 1:0] SAXIHP3BRESP,
    output logic        SAXIHP3BVALID,
    output logic [ 2:0] SAXIHP3RACOUNT,
    output logic [ 7:0] SAXIHP3RCOUNT,
    output logic [63:0] SAXIHP3RDATA,
    output logic [ 5:0] SAXIHP3RID,
    output logic        SAXIHP3RLAST,
    output logic [ 1:0] SAXIHP3RRESP,
    output logic        SAXIHP3RVALID,
    output logic [ 5:0] SAXIHP3WACOUNT,
    output logic [ 7:0] SAXIHP3WCOUNT,
    output logic        SAXIHP3WREADY,
    /* verilator lint_on UNDRIVEN */

    inout  logic [14:0] DDRA,
    inout  logic [ 2:0] DDRBA,
    inout  logic        DDRCASB,
    inout  logic        DDRCKE,
    inout  logic        DDRCKN,
    inout  logic        DDRCKP,
    inout  logic        DDRCSB,
    inout  logic [ 3:0] DDRDM,
    inout  logic [31:0] DDRDQ,
    inout  logic [ 3:0] DDRDQSN,
    inout  logic [ 3:0] DDRDQSP,
    inout  logic        DDRDRSTB,
    inout  logic        DDRODT,
    inout  logic        DDRRASB,
    inout  logic        DDRVRN,
    inout  logic        DDRVRP,
    inout  logic        DDRWEB,
    inout  logic [53:0] MIO,
    inout  logic        PSCLK,
    inout  logic        PSPORB,
    inout  logic        PSSRSTB,
    
    input  wire logic [ 3:0] DDRARB,
    input  wire logic        DMA0ACLK,
    input  wire logic        DMA0DAREADY,
    input  wire logic        DMA0DRLAST,
    input  wire logic [ 1:0] DMA0DRTYPE,
    input  wire logic        DMA0DRVALID,
    input  wire logic        DMA1ACLK,
    input  wire logic        DMA1DAREADY,
    input  wire logic        DMA1DRLAST,
    input  wire logic [ 1:0] DMA1DRTYPE,
    input  wire logic        DMA1DRVALID,
    input  wire logic        DMA2ACLK,
    input  wire logic        DMA2DAREADY,
    input  wire logic        DMA2DRLAST,
    input  wire logic [ 1:0] DMA2DRTYPE,
    input  wire logic        DMA2DRVALID,
    input  wire logic        DMA3ACLK,
    input  wire logic        DMA3DAREADY,
    input  wire logic        DMA3DRLAST,
    input  wire logic [ 1:0] DMA3DRTYPE,
    input  wire logic        DMA3DRVALID,
    input  wire logic        EMIOCAN0PHYRX,
    input  wire logic        EMIOCAN1PHYRX,
    input  wire logic        EMIOENET0EXTINTIN,
    input  wire logic        EMIOENET0GMIICOL,
    input  wire logic        EMIOENET0GMIICRS,
    input  wire logic        EMIOENET0GMIIRXCLK,
    input  wire logic [ 7:0] EMIOENET0GMIIRXD,
    input  wire logic        EMIOENET0GMIIRXDV,
    input  wire logic        EMIOENET0GMIIRXER,
    input  wire logic        EMIOENET0GMIITXCLK,
    input  wire logic        EMIOENET0MDIOI,
    input  wire logic        EMIOENET1EXTINTIN,
    input  wire logic        EMIOENET1GMIICOL,
    input  wire logic        EMIOENET1GMIICRS,
    input  wire logic        EMIOENET1GMIIRXCLK,
    input  wire logic [ 7:0] EMIOENET1GMIIRXD,
    input  wire logic        EMIOENET1GMIIRXDV,
    input  wire logic        EMIOENET1GMIIRXER,
    input  wire logic        EMIOENET1GMIITXCLK,
    input  wire logic        EMIOENET1MDIOI,
    input  wire logic [63:0] EMIOGPIOI,
    input  wire logic        EMIOI2C0SCLI,
    input  wire logic        EMIOI2C0SDAI,
    input  wire logic        EMIOI2C1SCLI,
    input  wire logic        EMIOI2C1SDAI,
    input  wire logic        EMIOPJTAGTCK,
    input  wire logic        EMIOPJTAGTDI,
    input  wire logic        EMIOPJTAGTMS,
    input  wire logic        EMIOSDIO0CDN,
    input  wire logic        EMIOSDIO0CLKFB,
    input  wire logic        EMIOSDIO0CMDI,
    input  wire logic [ 3:0] EMIOSDIO0DATAI,
    input  wire logic        EMIOSDIO0WP,
    input  wire logic        EMIOSDIO1CDN,
    input  wire logic        EMIOSDIO1CLKFB,
    input  wire logic        EMIOSDIO1CMDI,
    input  wire logic [ 3:0] EMIOSDIO1DATAI,
    input  wire logic        EMIOSDIO1WP,
    input  wire logic        EMIOSPI0MI,
    input  wire logic        EMIOSPI0SCLKI,
    input  wire logic        EMIOSPI0SI,
    input  wire logic        EMIOSPI0SSIN,
    input  wire logic        EMIOSPI1MI,
    input  wire logic        EMIOSPI1SCLKI,
    input  wire logic        EMIOSPI1SI,
    input  wire logic        EMIOSPI1SSIN,
    input  wire logic        EMIOSRAMINTIN,
    input  wire logic        EMIOTRACECLK,
    input  wire logic [ 2:0] EMIOTTC0CLKI,
    input  wire logic [ 2:0] EMIOTTC1CLKI,
    input  wire logic        EMIOUART0CTSN,
    input  wire logic        EMIOUART0DCDN,
    input  wire logic        EMIOUART0DSRN,
    input  wire logic        EMIOUART0RIN,
    input  wire logic        EMIOUART0RX,
    input  wire logic        EMIOUART1CTSN,
    input  wire logic        EMIOUART1DCDN,
    input  wire logic        EMIOUART1DSRN,
    input  wire logic        EMIOUART1RIN,
    input  wire logic        EMIOUART1RX,
    input  wire logic        EMIOUSB0VBUSPWRFAULT,
    input  wire logic        EMIOUSB1VBUSPWRFAULT,
    input  wire logic        EMIOWDTCLKI,
    input  wire logic        EVENTEVENTI,
    input  wire logic [ 3:0] FCLKCLKTRIGN,
    input  wire logic        FPGAIDLEN,
    input  wire logic [ 3:0] FTMDTRACEINATID,
    input  wire logic        FTMDTRACEINCLOCK,
    input  wire logic [31:0] FTMDTRACEINDATA,
    input  wire logic        FTMDTRACEINVALID,
    input  wire logic [31:0] FTMTF2PDEBUG,
    input  wire logic [ 3:0] FTMTF2PTRIG,
    input  wire logic [ 3:0] FTMTP2FTRIGACK,
    input  wire logic [19:0] IRQF2P,
    input  wire logic        MAXIGP0ACLK,
    input  wire logic        MAXIGP0ARREADY,
    input  wire logic        MAXIGP0AWREADY,
    input  wire logic [11:0] MAXIGP0BID,
    input  wire logic [ 1:0] MAXIGP0BRESP,
    input  wire logic        MAXIGP0BVALID,
    input  wire logic [31:0] MAXIGP0RDATA,
    input  wire logic [11:0] MAXIGP0RID,
    input  wire logic        MAXIGP0RLAST,
    input  wire logic [ 1:0] MAXIGP0RRESP,
    input  wire logic        MAXIGP0RVALID,
    input  wire logic        MAXIGP0WREADY,
    input  wire logic        MAXIGP1ACLK,
    input  wire logic        MAXIGP1ARREADY,
    input  wire logic        MAXIGP1AWREADY,
    input  wire logic [11:0] MAXIGP1BID,
    input  wire logic [ 1:0] MAXIGP1BRESP,
    input  wire logic        MAXIGP1BVALID,
    input  wire logic [31:0] MAXIGP1RDATA,
    input  wire logic [11:0] MAXIGP1RID,
    input  wire logic        MAXIGP1RLAST,
    input  wire logic [ 1:0] MAXIGP1RRESP,
    input  wire logic        MAXIGP1RVALID,
    input  wire logic        MAXIGP1WREADY,
    input  wire logic        SAXIACPACLK,
    input  wire logic [31:0] SAXIACPARADDR,
    input  wire logic [ 1:0] SAXIACPARBURST,
    input  wire logic [ 3:0] SAXIACPARCACHE,
    input  wire logic [ 2:0] SAXIACPARID,
    input  wire logic [ 3:0] SAXIACPARLEN,
    input  wire logic [ 1:0] SAXIACPARLOCK,
    input  wire logic [ 2:0] SAXIACPARPROT,
    input  wire logic [ 3:0] SAXIACPARQOS,
    input  wire logic [ 1:0] SAXIACPARSIZE,
    input  wire logic [ 4:0] SAXIACPARUSER,
    input  wire logic        SAXIACPARVALID,
    input  wire logic [31:0] SAXIACPAWADDR,
    input  wire logic [ 1:0] SAXIACPAWBURST,
    input  wire logic [ 3:0] SAXIACPAWCACHE,
    input  wire logic [ 2:0] SAXIACPAWID,
    input  wire logic [ 3:0] SAXIACPAWLEN,
    input  wire logic [ 1:0] SAXIACPAWLOCK,
    input  wire logic [ 2:0] SAXIACPAWPROT,
    input  wire logic [ 3:0] SAXIACPAWQOS,
    input  wire logic [ 1:0] SAXIACPAWSIZE,
    input  wire logic [ 4:0] SAXIACPAWUSER,
    input  wire logic        SAXIACPAWVALID,
    input  wire logic        SAXIACPBREADY,
    input  wire logic        SAXIACPRREADY,
    input  wire logic [63:0] SAXIACPWDATA,
    input  wire logic [ 2:0] SAXIACPWID,
    input  wire logic        SAXIACPWLAST,
    input  wire logic [ 7:0] SAXIACPWSTRB,
    input  wire logic        SAXIACPWVALID,
    input  wire logic        SAXIGP0ACLK,
    input  wire logic [31:0] SAXIGP0ARADDR,
    input  wire logic [ 1:0] SAXIGP0ARBURST,
    input  wire logic [ 3:0] SAXIGP0ARCACHE,
    input  wire logic [ 5:0] SAXIGP0ARID,
    input  wire logic [ 3:0] SAXIGP0ARLEN,
    input  wire logic [ 1:0] SAXIGP0ARLOCK,
    input  wire logic [ 2:0] SAXIGP0ARPROT,
    input  wire logic [ 3:0] SAXIGP0ARQOS,
    input  wire logic [ 1:0] SAXIGP0ARSIZE,
    input  wire logic        SAXIGP0ARVALID,
    input  wire logic [31:0] SAXIGP0AWADDR,
    input  wire logic [ 1:0] SAXIGP0AWBURST,
    input  wire logic [ 3:0] SAXIGP0AWCACHE,
    input  wire logic [ 5:0] SAXIGP0AWID,
    input  wire logic [ 3:0] SAXIGP0AWLEN,
    input  wire logic [ 1:0] SAXIGP0AWLOCK,
    input  wire logic [ 2:0] SAXIGP0AWPROT,
    input  wire logic [ 3:0] SAXIGP0AWQOS,
    input  wire logic [ 1:0] SAXIGP0AWSIZE,
    input  wire logic        SAXIGP0AWVALID,
    input  wire logic        SAXIGP0BREADY,
    input  wire logic        SAXIGP0RREADY,
    input  wire logic [31:0] SAXIGP0WDATA,
    input  wire logic [ 5:0] SAXIGP0WID,
    input  wire logic        SAXIGP0WLAST,
    input  wire logic [ 3:0] SAXIGP0WSTRB,
    input  wire logic        SAXIGP0WVALID,
    input  wire logic        SAXIGP1ACLK,
    input  wire logic [31:0] SAXIGP1ARADDR,
    input  wire logic [ 1:0] SAXIGP1ARBURST,
    input  wire logic [ 3:0] SAXIGP1ARCACHE,
    input  wire logic [ 5:0] SAXIGP1ARID,
    input  wire logic [ 3:0] SAXIGP1ARLEN,
    input  wire logic [ 1:0] SAXIGP1ARLOCK,
    input  wire logic [ 2:0] SAXIGP1ARPROT,
    input  wire logic [ 3:0] SAXIGP1ARQOS,
    input  wire logic [ 1:0] SAXIGP1ARSIZE,
    input  wire logic        SAXIGP1ARVALID,
    input  wire logic [31:0] SAXIGP1AWADDR,
    input  wire logic [ 1:0] SAXIGP1AWBURST,
    input  wire logic [ 3:0] SAXIGP1AWCACHE,
    input  wire logic [ 5:0] SAXIGP1AWID,
    input  wire logic [ 3:0] SAXIGP1AWLEN,
    input  wire logic [ 1:0] SAXIGP1AWLOCK,
    input  wire logic [ 2:0] SAXIGP1AWPROT,
    input  wire logic [ 3:0] SAXIGP1AWQOS,
    input  wire logic [ 1:0] SAXIGP1AWSIZE,
    input  wire logic        SAXIGP1AWVALID,
    input  wire logic        SAXIGP1BREADY,
    input  wire logic        SAXIGP1RREADY,
    input  wire logic [31:0] SAXIGP1WDATA,
    input  wire logic [ 5:0] SAXIGP1WID,
    input  wire logic        SAXIGP1WLAST,
    input  wire logic [ 3:0] SAXIGP1WSTRB,
    input  wire logic        SAXIGP1WVALID,
    input  wire logic        SAXIHP0ACLK,
    input  wire logic [31:0] SAXIHP0ARADDR,
    input  wire logic [ 1:0] SAXIHP0ARBURST,
    input  wire logic [ 3:0] SAXIHP0ARCACHE,
    input  wire logic [ 5:0] SAXIHP0ARID,
    input  wire logic [ 3:0] SAXIHP0ARLEN,
    input  wire logic [ 1:0] SAXIHP0ARLOCK,
    input  wire logic [ 2:0] SAXIHP0ARPROT,
    input  wire logic [ 3:0] SAXIHP0ARQOS,
    input  wire logic [ 1:0] SAXIHP0ARSIZE,
    input  wire logic        SAXIHP0ARVALID,
    input  wire logic [31:0] SAXIHP0AWADDR,
    input  wire logic [ 1:0] SAXIHP0AWBURST,
    input  wire logic [ 3:0] SAXIHP0AWCACHE,
    input  wire logic [ 5:0] SAXIHP0AWID,
    input  wire logic [ 3:0] SAXIHP0AWLEN,
    input  wire logic [ 1:0] SAXIHP0AWLOCK,
    input  wire logic [ 2:0] SAXIHP0AWPROT,
    input  wire logic [ 3:0] SAXIHP0AWQOS,
    input  wire logic [ 1:0] SAXIHP0AWSIZE,
    input  wire logic        SAXIHP0AWVALID,
    input  wire logic        SAXIHP0BREADY,
    input  wire logic        SAXIHP0RDISSUECAP1EN,
    input  wire logic        SAXIHP0RREADY,
    input  wire logic [63:0] SAXIHP0WDATA,
    input  wire logic [ 5:0] SAXIHP0WID,
    input  wire logic        SAXIHP0WLAST,
    input  wire logic        SAXIHP0WRISSUECAP1EN,
    input  wire logic [ 7:0] SAXIHP0WSTRB,
    input  wire logic        SAXIHP0WVALID,
    input  wire logic        SAXIHP1ACLK,
    input  wire logic [31:0] SAXIHP1ARADDR,
    input  wire logic [ 1:0] SAXIHP1ARBURST,
    input  wire logic [ 3:0] SAXIHP1ARCACHE,
    input  wire logic [ 5:0] SAXIHP1ARID,
    input  wire logic [ 3:0] SAXIHP1ARLEN,
    input  wire logic [ 1:0] SAXIHP1ARLOCK,
    input  wire logic [ 2:0] SAXIHP1ARPROT,
    input  wire logic [ 3:0] SAXIHP1ARQOS,
    input  wire logic [ 1:0] SAXIHP1ARSIZE,
    input  wire logic        SAXIHP1ARVALID,
    input  wire logic [31:0] SAXIHP1AWADDR,
    input  wire logic [ 1:0] SAXIHP1AWBURST,
    input  wire logic [ 3:0] SAXIHP1AWCACHE,
    input  wire logic [ 5:0] SAXIHP1AWID,
    input  wire logic [ 3:0] SAXIHP1AWLEN,
    input  wire logic [ 1:0] SAXIHP1AWLOCK,
    input  wire logic [ 2:0] SAXIHP1AWPROT,
    input  wire logic [ 3:0] SAXIHP1AWQOS,
    input  wire logic [ 1:0] SAXIHP1AWSIZE,
    input  wire logic        SAXIHP1AWVALID,
    input  wire logic        SAXIHP1BREADY,
    input  wire logic        SAXIHP1RDISSUECAP1EN,
    input  wire logic        SAXIHP1RREADY,
    input  wire logic [63:0] SAXIHP1WDATA,
    input  wire logic [ 5:0] SAXIHP1WID,
    input  wire logic        SAXIHP1WLAST,
    input  wire logic        SAXIHP1WRISSUECAP1EN,
    input  wire logic [ 7:0] SAXIHP1WSTRB,
    input  wire logic        SAXIHP1WVALID,
    input  wire logic        SAXIHP2ACLK,
    input  wire logic [31:0] SAXIHP2ARADDR,
    input  wire logic [ 1:0] SAXIHP2ARBURST,
    input  wire logic [ 3:0] SAXIHP2ARCACHE,
    input  wire logic [ 5:0] SAXIHP2ARID,
    input  wire logic [ 3:0] SAXIHP2ARLEN,
    input  wire logic [ 1:0] SAXIHP2ARLOCK,
    input  wire logic [ 2:0] SAXIHP2ARPROT,
    input  wire logic [ 3:0] SAXIHP2ARQOS,
    input  wire logic [ 1:0] SAXIHP2ARSIZE,
    input  wire logic        SAXIHP2ARVALID,
    input  wire logic [31:0] SAXIHP2AWADDR,
    input  wire logic [ 1:0] SAXIHP2AWBURST,
    input  wire logic [ 3:0] SAXIHP2AWCACHE,
    input  wire logic [ 5:0] SAXIHP2AWID,
    input  wire logic [ 3:0] SAXIHP2AWLEN,
    input  wire logic [ 1:0] SAXIHP2AWLOCK,
    input  wire logic [ 2:0] SAXIHP2AWPROT,
    input  wire logic [ 3:0] SAXIHP2AWQOS,
    input  wire logic [ 1:0] SAXIHP2AWSIZE,
    input  wire logic        SAXIHP2AWVALID,
    input  wire logic        SAXIHP2BREADY,
    input  wire logic        SAXIHP2RDISSUECAP1EN,
    input  wire logic        SAXIHP2RREADY,
    input  wire logic [63:0] SAXIHP2WDATA,
    input  wire logic [ 5:0] SAXIHP2WID,
    input  wire logic        SAXIHP2WLAST,
    input  wire logic        SAXIHP2WRISSUECAP1EN,
    input  wire logic [ 7:0] SAXIHP2WSTRB,
    input  wire logic        SAXIHP2WVALID,
    input  wire logic        SAXIHP3ACLK,
    input  wire logic [31:0] SAXIHP3ARADDR,
    input  wire logic [ 1:0] SAXIHP3ARBURST,
    input  wire logic [ 3:0] SAXIHP3ARCACHE,
    input  wire logic [ 5:0] SAXIHP3ARID,
    input  wire logic [ 3:0] SAXIHP3ARLEN,
    input  wire logic [ 1:0] SAXIHP3ARLOCK,
    input  wire logic [ 2:0] SAXIHP3ARPROT,
    input  wire logic [ 3:0] SAXIHP3ARQOS,
    input  wire logic [ 1:0] SAXIHP3ARSIZE,
    input  wire logic        SAXIHP3ARVALID,
    input  wire logic [31:0] SAXIHP3AWADDR,
    input  wire logic [ 1:0] SAXIHP3AWBURST,
    input  wire logic [ 3:0] SAXIHP3AWCACHE,
    input  wire logic [ 5:0] SAXIHP3AWID,
    input  wire logic [ 3:0] SAXIHP3AWLEN,
    input  wire logic [ 1:0] SAXIHP3AWLOCK,
    input  wire logic [ 2:0] SAXIHP3AWPROT,
    input  wire logic [ 3:0] SAXIHP3AWQOS,
    input  wire logic [ 1:0] SAXIHP3AWSIZE,
    input  wire logic        SAXIHP3AWVALID,
    input  wire logic        SAXIHP3BREADY,
    input  wire logic        SAXIHP3RDISSUECAP1EN,
    input  wire logic        SAXIHP3RREADY,
    input  wire logic [63:0] SAXIHP3WDATA,
    input  wire logic [ 5:0] SAXIHP3WID,
    input  wire logic        SAXIHP3WLAST,
    input  wire logic        SAXIHP3WRISSUECAP1EN,
    input  wire logic [ 7:0] SAXIHP3WSTRB,
    input  wire logic        SAXIHP3WVALID
    /* verilator lint_on UNUSED */
);

    // Null module

endmodule
