//
//    Copyright (C) 2022  Jakub Hladik
//
//    This program is free software: you can redistribute it and/or modify
//    it under the terms of the GNU General Public License as published by
//    the Free Software Foundation, either version 3 of the License, or
//    (at your option) any later version.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    You should have received a copy of the GNU General Public License
//    along with this program.  If not, see <https://www.gnu.org/licenses/>.
//

`default_nettype none

module OBUFDS #(
    /* verilator lint_off UNUSED */
    parameter IOSTANDARD = "DEFAULT",
    parameter SLEW       = "SLOW"
    /* verilator lint_on UNUSED */
) (
    /* verilator lint_off UNUSED */
    /* verilator lint_off UNDRIVEN */
    output      logic O,
    output      logic OB,
    /* verilator lint_on UNDRIVEN */
    input  wire logic I
    /* verilator lint_on UNUSED */
);

    // Null module

endmodule
